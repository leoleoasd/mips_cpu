module mips(
    input clk,
    input rst
);

endmodule